package lns_mac_pkg;


parameter IN_BITS = 15; 
parameter OUT_BITS = 15;
parameter NUM_DATA_IN = 32;

endpackage
